module encoder_8(d,a,b,c);
input [7:0]d;
output a,b,c;



endmodule
