module mux_8(s0,s1,s2,d,y);
input s0,s1,s2;
input [7:0]d;
output y;



endmodule
