module decoder_8(a,b,c,y);
input a,b,c;
output[7:0]y;



endmodule
