module demux_8(s,d,y);
input [2:0]s;
input d;
output [7:0]y;




endmodule
